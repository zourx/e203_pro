 /*                                                                      
 Copyright 2018 Nuclei System Technology, Inc.                
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
  Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */                                                                      
                                                                         
                                                                         
                                                                         
//=====================================================================
//
// Designer   : Bob Hu
//
// Description:
//  The top level module of plic
//
// ====================================================================

`include "e203_defines.v"

module sirv_plic_top(
  input   clk,
  input   rst_n,

  input                      i_icb_cmd_valid,
  output                     i_icb_cmd_ready,
  input  [32-1:0]            i_icb_cmd_addr, 
  input                      i_icb_cmd_read, 
  input  [32-1:0]            i_icb_cmd_wdata,
  
  output                     i_icb_rsp_valid,
  input                      i_icb_rsp_ready,
  output [32-1:0]            i_icb_rsp_rdata,

  input   io_devices_0_0,
  input   io_devices_0_1,
  input   io_devices_0_2,
  input   io_devices_0_3,
  input   io_devices_0_4,
  input   io_devices_0_5,
  input   io_devices_0_6,
  input   io_devices_0_7,
  input   io_devices_0_8,
  input   io_devices_0_9,
  input   io_devices_0_10,
  input   io_devices_0_11,
  input   io_devices_0_12,
  input   io_devices_0_13,
  input   io_devices_0_14,
  input   io_devices_0_15,
  input   io_devices_0_16,
  input   io_devices_0_17,
  input   io_devices_0_18,
  input   io_devices_0_19,
  input   io_devices_0_20,
  input   io_devices_0_21,
  input   io_devices_0_22,
  input   io_devices_0_23,
  input   io_devices_0_24,
  input   io_devices_0_25,
  input   io_devices_0_26,
  input   io_devices_0_27,
  input   io_devices_0_28,
  input   io_devices_0_29,
  input   io_devices_0_30,
  input   io_devices_0_31,
  input   io_devices_0_32,
  input   io_devices_0_33,
  input   io_devices_0_34,
  input   io_devices_0_35,
  input   io_devices_0_36,
  input   io_devices_0_37,
  input   io_devices_0_38,
  input   io_devices_0_39,
  input   io_devices_0_40,
  input   io_devices_0_41,
  input   io_devices_0_42,
  input   io_devices_0_43,
  input   io_devices_0_44,
  input   io_devices_0_45,
  input   io_devices_0_46,
  input   io_devices_0_47,
  input   io_devices_0_48,
  input   io_devices_0_49,
  input   io_devices_0_50,
  input   io_devices_0_51,
  output  io_harts_0_0,

/// nts
  input        saveregdone_2nplic,
  output [2:0] iq_aftrap_nplic2nts,
  input  [1:0] trap_stage_nts2nplic,
  output [1:0] trap_type2core,

/// to nplic
  input                  ret2nplic,
  input [3:0]            num_trap2nplic,
  input                  nts_full_o2nplic,
  input [`E203_XLEN-1:0] x2_sp,

  output bftail_trap,
  output nest_trap_2ntsctrl,
  input  aftail_trap,

/// clint
  input                          tm_stop,

  input                          clint_icb_cmd_valid,
  output                         clint_icb_cmd_ready,
  input  [`E203_ADDR_SIZE-1:0]   clint_icb_cmd_addr, 
  input                          clint_icb_cmd_read, 
  input  [`E203_XLEN-1:0]        clint_icb_cmd_wdata,
  input  [`E203_XLEN/8-1:0]      clint_icb_cmd_wmask,

  output                         clint_icb_rsp_valid,
  input                          clint_icb_rsp_ready,
  output                         clint_icb_rsp_err,
  output [`E203_XLEN-1:0]        clint_icb_rsp_rdata,

  output                         clint_tmr_irq,
  output                         clint_sft_irq,

  input                          aon_rtcToggle_a,
  input [31:0]                   console_icb_cmd_wdata 

);


///////////////////////////////////////////////////////////////////////////////////////////////////////////////
/// nts test
  reg [31:0] count;
  always @(posedge clk or negedge rst_n) begin
    if (~rst_n) begin
      count <= 'd0;
    end if (count < 'h499999) begin
      count <= count + 1'd1;
    end else begin
      count <= 'b0;
    end
  end

  assign plic_irq_i         = (plic_irq_i_device != 0) ? interrupt_test_irq : plic_irq_i_device;
  assign io_harts_0_0       = plic_irq;

  wire                    plic_irq;
  wire [PLIC_IRQ_NUM-1:0] plic_irq_i;
  wire [PLIC_IRQ_NUM-1:0] interrupt_test_irq;
  wire                    interrupt_test;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// 追咬尾 T -> E -> T
// platfrom.h
// #define CLINT_TIMEBASE_FREQ 10000



  // assign interrupt_test     = ((count == 32'd91618)) ? 1'b1 : 1'b0;

  // assign interrupt_test_irq = (interrupt_test & (count == 32'd91618)) ? (53'h1 << 14) :  53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// 巢狀 T -> E
// platfrom.h
// #define CLINT_TIMEBASE_FREQ 10000



  // assign interrupt_test     = ((count == 32'd91690)) ? 1'b1 : 1'b0;

  // assign interrupt_test_irq = (interrupt_test & (count == 32'd91690)) ? (53'h1 << 14) :  53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// 巢狀 S -> E
// sched.c - cls task_yield
// void user_task1(void)
// { task_yield(); }

// user.c  - op  MSIP = 1
// void task_yield()
// { *(uint32_t*)CLINT_MSIP(id) = 1;}



  // assign interrupt_test     = ((count == 32'd83540)) ? 1'b1 : 1'b0;

  // assign interrupt_test_irq = (interrupt_test & (count == 32'd83540)) ? (53'h1 << 14) :  53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// 追咬尾 S -> E -> S
// sched.c - cls task_yield
// void user_task1(void)
// { task_yield(); }

// user.c  - op  MSIP = 1
// void task_yield()
// { *(uint32_t*)CLINT_MSIP(id) = 1;}



  // assign interrupt_test     = ((count == 32'd83524)) ? 1'b1 : 1'b0;

  // assign interrupt_test_irq = (interrupt_test & (count == 32'd83524)) ? (53'h1 << 14) :  53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// E -> E -> E

  // assign interrupt_test     = ((count == 32'd83460)
  //                             |(count == 32'd83463)) ? 1'b1 : 1'b0;

  // assign interrupt_test_irq = (interrupt_test & (count == 32'd83460)) ? (53'h1 << 14) : 
  //                             (interrupt_test & (count == 32'd83463)) ? (53'h1 << 13) :  53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////
//// 巢狀 full

  assign interrupt_test     = ((count == 32'd98819)
                              |(count == 32'd98849)
                              |(count == 32'd98879)
                              |(count == 32'd98909)
                              |(count == 32'd98939)
                              |(count == 32'd98969)
                              |(count == 32'd98999)
                              |(count == 32'd99029)
                              |(count == 32'd99059)
                              |(count == 32'd99079)
                              |(count == 32'd99109)
                              |(count == 32'd99139)
                              |(count == 32'd99149)) ? 1'b1 : 1'b0;

  assign interrupt_test_irq = (interrupt_test & (count == 32'd98819)) ? (53'h1 << 14) :
                              (interrupt_test & (count == 32'd98849)) ? (53'h1 << 13) : 
                              (interrupt_test & (count == 32'd98879)) ? (53'h1 << 12) :
                              (interrupt_test & (count == 32'd98909)) ? (53'h1 << 11) : 
                              (interrupt_test & (count == 32'd98939)) ? (53'h1 << 10) : 
                              (interrupt_test & (count == 32'd98969)) ? (53'h1 <<  9) :
                              (interrupt_test & (count == 32'd98999)) ? (53'h1 <<  8) : 
                              (interrupt_test & (count == 32'd99029)) ? (53'h1 <<  7) : 
                              (interrupt_test & (count == 32'd99059)) ? (53'h1 <<  6) :
                              (interrupt_test & (count == 32'd99079)) ? (53'h1 <<  5) : 
                              (interrupt_test & (count == 32'd99109)) ? (53'h1 <<  4) : 
                              (interrupt_test & (count == 32'd99139)) ? (53'h1 <<  3) :
                              (interrupt_test & (count == 32'd99149)) ? (53'h1 <<  2) : 53'h0;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////


localparam PLIC_IRQ_NUM = 53;// The number can be enlarged as long as not larger than 1024
wire [PLIC_IRQ_NUM-1:0] plic_irq_i_device = { 
                  io_devices_0_51  ,
                  io_devices_0_50  ,

                  io_devices_0_49  ,
                  io_devices_0_48  ,
                  io_devices_0_47  ,
                  io_devices_0_46  ,
                  io_devices_0_45  ,
                  io_devices_0_44  ,
                  io_devices_0_43  ,
                  io_devices_0_42  ,
                  io_devices_0_41  ,
                  io_devices_0_40  ,

                  io_devices_0_39  ,
                  io_devices_0_38  ,
                  io_devices_0_37  ,
                  io_devices_0_36  ,
                  io_devices_0_35  ,
                  io_devices_0_34  ,
                  io_devices_0_33  ,
                  io_devices_0_32  ,
                  io_devices_0_31  ,
                  io_devices_0_30  ,

                  io_devices_0_29  ,
                  io_devices_0_28  ,
                  io_devices_0_27  ,
                  io_devices_0_26  ,
                  io_devices_0_25  ,
                  io_devices_0_24  ,
                  io_devices_0_23  ,
                  io_devices_0_22  ,
                  io_devices_0_21  ,
                  io_devices_0_20  ,

                  io_devices_0_19  ,
                  io_devices_0_18  ,
                  io_devices_0_17  ,
                  io_devices_0_16  ,
                  io_devices_0_15  ,
                  io_devices_0_14  ,
                  io_devices_0_13  ,
                  io_devices_0_12  ,
                  io_devices_0_11  ,
                  io_devices_0_10  ,

                  io_devices_0_9  ,
                  io_devices_0_8  ,
                  io_devices_0_7  ,
                  io_devices_0_6  ,
                  io_devices_0_5  ,
                  io_devices_0_4  ,
                  io_devices_0_3  ,
                  io_devices_0_2  ,
                  io_devices_0_1  ,
                  io_devices_0_0  ,

                  1'b0 };// The IRQ0 must be tied to zero

wire [31:0] plic_addr = (i_icb_cmd_addr[31:24] == 'b00010001) ? 'b0 : i_icb_cmd_addr; 

sirv_plic_man #(
    .PLIC_PRIO_WIDTH   (3),
    .PLIC_IRQ_NUM      (PLIC_IRQ_NUM),
    .PLIC_IRQ_NUM_LOG2 (6),
    .PLIC_ICB_RSP_FLOP (1),
    .PLIC_IRQ_I_FLOP   (1),
    .PLIC_IRQ_O_FLOP   (1) 
) u_sirv_plic_man(
    .clk              (clk            ),      
    .rst_n            (rst_n          ),

    .icb_cmd_valid  (i_icb_cmd_valid),
    .icb_cmd_addr   (plic_addr[24-1:0] ),
    .icb_cmd_read   (i_icb_cmd_read ),
    .icb_cmd_wdata  (i_icb_cmd_wdata),
    .icb_rsp_ready  (i_icb_rsp_ready),
                    
    .icb_rsp_valid  (i_icb_rsp_valid),
    .icb_cmd_ready  (i_icb_cmd_ready),
    .icb_rsp_rdata  (i_icb_rsp_rdata),

    .plic_irq_i (plic_irq_i),
    .plic_irq_o (plic_irq   ),

/// nts
    .bftail_trap          (bftail_trap          ),
    .nest_trap_2ntsctrl   (nest_trap_2ntsctrl   ),
    .aftail_trap          (aftail_trap          ),
    .iq_aftrap_nplic2nts  (iq_aftrap_nplic2nts  ),
    .saveregdone_2nplic   (saveregdone_2nplic   ),
    .trap_stage_nts2nplic (trap_stage_nts2nplic ),
    .trap_type2core       (trap_type2core       ),

/// to nplic
    .ret2nplic            (ret2nplic),
    .num_trap2nplic       (num_trap2nplic),
    .nts_full_o2nplic     (nts_full_o2nplic),
    .x2_sp                (x2_sp),

/// clint
    .tm_stop              (tm_stop),

    .clint_icb_cmd_valid  (clint_icb_cmd_valid),
    .clint_icb_cmd_ready  (clint_icb_cmd_ready),
    .clint_icb_cmd_addr   (clint_icb_cmd_addr ),
    .clint_icb_cmd_read   (clint_icb_cmd_read ),
    .clint_icb_cmd_wdata  (clint_icb_cmd_wdata),
    .clint_icb_cmd_wmask  (clint_icb_cmd_wmask),
    
    .clint_icb_rsp_valid  (clint_icb_rsp_valid),
    .clint_icb_rsp_ready  (clint_icb_rsp_ready),
    .clint_icb_rsp_err    (clint_icb_rsp_err  ),
    .clint_icb_rsp_rdata  (clint_icb_rsp_rdata),

    .clint_tmr_irq        (clint_tmr_irq),
    .clint_sft_irq        (clint_sft_irq),

    .aon_rtcToggle_a      (aon_rtcToggle_a)
);

endmodule
